module and2
(
    input wire [1:0]in0,
    input wire [1:0] in1,
    output wire [1:0] out
);
  assign  out=in0&in1;
endmodule